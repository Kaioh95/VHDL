library ieee;
use ieee.std_logic_1164.all;

entity demux_1x4_ite is 
	port(
		a: in std_logic;
		s0, s1: in std_logic;
		o0, o1, o2, o3: out std_logic
	);

end demux_1x4_ite;

architecture arch of demux_1x4_ite is
	begin
		process (a, s0, s1) is
		begin
			if(s1='0' and s0='0') then
				o0 <= '1';
				o1 <= '0';
				o2 <= '0';
				o3 <= '0';
			elsif(s1='0' and s0='1') then
				o0 <= '0';
				o1 <= '1';
				o2 <= '0';
				o3 <= '0';
			elsif(s1='1' and s0='0') then
				o0 <= '0';
				o1 <= '0';
				o2 <= '1';
				o3 <= '0';
			elsif(s1='1' and s0='1') then
				o0 <= '0';
				o1 <= '0';
				o2 <= '0';
				o3 <= '1';
			end if;
		end process;
	end arch;